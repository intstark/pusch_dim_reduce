module pus_rst (
		output wire [15:0] source,     //    sources.source
		input  wire        source_clk  // source_clk.clk
	);
endmodule

