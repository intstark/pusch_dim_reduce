// rom_65536x64_L0.v

// Generated using ACDS version 23.2 94

`timescale 1 ps / 1 ps
module rom_65536x64_L0 (
		output wire [63:0] q,       //       q.dataout
		input  wire [15:0] address, // address.address
		input  wire        clock,   //   clock.clk
		input  wire        rden     //    rden.rden
	);

	rom_65536x64_L0_rom_1port_2020_opruxui rom_1port_0 (
		.q       (q),       //  output,  width = 64,       q.dataout
		.address (address), //   input,  width = 16, address.address
		.clock   (clock),   //   input,   width = 1,   clock.clk
		.rden    (rden)     //   input,   width = 1,    rden.rden
	);

endmodule
